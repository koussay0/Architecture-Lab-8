
`timescale 1ns / 1ps

module InstMem (input [5:0] offset, output [31:0] data_out);

   //Instruction Memory
   reg [31:0] mem [0:63];
   assign data_out = mem[offset];
   initial begin
//    mem[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0,
//    mem[1]=32'b00000000000000000010000010000011 ; //lw x1, 0(x0) x1= 17
//    mem[2]=32'b00000000000000000000000000110011 ; //add x0, x0, x0
//    mem[3]=32'b00000000000000000000000000110011 ; //add x0, x0, x0 
//    mem[4]=32'b00000000000000000000000000110011 ; //add x0, x0, x0 
//    mem[5]=32'b00000000010000000010000100000011 ; //lw x2, 4(x0)  x2 = 9 
//    mem[6]=32'b00000000000000000000000000110011 ; //add x0, x0, x0 
//    mem[7]=32'b00000000000000000000000000110011 ; //add x0, x0, x0
//    mem[8]=32'b00000000000000000000000000110011 ; //add x0, x0, x0 
//    mem[9]=32'b00000000100000000010000110000011 ; //lw x3, 8(x0) x3 = 25
//    mem[10]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[11]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[12]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[13]=32'b00000000001000001110001000110011 ; //or x4, x1, x2  x4 = 25 
//    mem[14]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[15]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[16]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[17]=32'b00000010001100100000000001100011; //beq x4, x3, 16 should branch 
//    mem[18]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[19]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[20]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[21]=32'b00000000001000001000000110110011 ; //add x3, x1, x2  x3 = 26 
//    mem[22]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[23]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[24]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[25]=32'b00000000001000011000001010110011 ; //add x5, x3, x2  x5 = 34 
//    mem[26]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[27]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[28]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[29]=32'b00000000010100000010011000100011; //sw x5, 12(x0)
//    mem[30]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[31]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[32]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//    mem[33]=32'b00000000110000000010001100000011 ; //lw x6, 12(x0)
//    mem[34]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[35]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[36]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[37]=32'b00000000000100110111001110110011 ; //and x7, x6, x1 
//    mem[38]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[39]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[40]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[41]=32'b01000000001000001000010000110011 ; //sub x8, x1, x2 
//    mem[42]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[43]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[44]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[45]=32'b00000000001000001000000000110011 ; //add x0, x1, x2 
//    mem[46]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[47]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[48]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
//    mem[49]=32'b00000000000100000000010010110011 ; //add x9, x0, x1end


    mem[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0,
    mem[1]=32'b00000000000000000010000010000011 ; //lw x1, 0(x0) x1= 17
    mem[2]=32'b00000000010000000010000100000011 ; //lw x2, 4(x0)  x2 = 9 
    mem[3]=32'b00000000100000000010000110000011 ; //lw x3, 8(x0) x3 = 25
    mem[4]=32'b00000000001000001110001000110011 ; //or x4, x1, x2  x4 = 25 
    mem[5]=32'b00000010001100100000000001100011; //beq x4, x3, 16 should branch 
    mem[6]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
    mem[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
    mem[8]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
    mem[9]=32'b00000000001000001000000110110011 ; //add x3, x1, x2  x3 = 26 
    mem[10]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
    mem[11]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
    mem[12]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
    mem[13]=32'b00000000001000011000001010110011 ; //add x5, x3, x2  x5 = 34 
    mem[14]=32'b00000000010100000010011000100011; //sw x5, 12(x0)
    mem[15]=32'b00000000110000000010001100000011 ; //lw x6, 12(x0)  34
     mem[16]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
    mem[17]=32'b00000000000100110111001110110011 ; //and x7, x6, x1 
    mem[18]=32'b01000000001000001000010000110011 ; //sub x8, x1, x2 
    mem[19]=32'b00000000000100000000010010110011 ; //add x9, x0, x1 end
   
  
    
    end
    
endmodule